// This is a minimal verilog module

module top;

endmodule

