/*
********************************************
* MODULE ice40_loopback.v
*
* This project is a test of the uart.
* It reads a character from the rx side
* of the uart then sends it on the tx side.
*
* Target Board: ICE40HX8K Breakout Board
*
* Author: Brandon Blodget
* Create Date: 06/09/2019
*
********************************************
*/

// Force error when implicit net has no type.
`default_nettype none

module ice40_loopback #
(
    parameter integer CLK_FREQUENCY = 96_000_000,
    parameter integer BAUD = 115_200,
    parameter integer NUM_LEDS = 8
)
(
    input wire  clk_12mhz,
    input wire reset_n,

    input wire  rxd,  // rxd
    output wire txd,  // txd

    output reg [7:0] led

);

/*
********************************************
* Signals
********************************************
*/

wire clk_96mhz;
wire locked;
wire reset;

reg uart_rd;
reg uart_wr;
wire rx_valid;
wire tx_busy;
reg [7:0] tx_data;
wire [7:0] rx_data;

/*
****************************
* Instantiations
****************************
*/

// Use PLL to get 50mhz clock
pll_96mhz pll_96mhz_inst (
    .clock_in(clk_12mhz),
    .clock_out(clk_96mhz),
    .locked(locked)
);

buart # (
    .CLKFREQ(CLK_FREQUENCY)
) uart_inst (
   .clk(clk_96mhz),
   .resetq(~reset),
   .baud(BAUD),
   .rx(rxd),           // recv wire
   .tx(txd),          // xmit wire
   .rd(uart_rd),           // read strobe
   .wr(uart_wr),           // write strobe
   .valid(rx_valid),       // has recv data 
   .busy(tx_busy),        // is transmitting
   .tx_data(tx_data),
   .rx_data(rx_data) // data
);

/*
****************************
* Main
****************************
*/

// Hold reset on power up then release.
// ice40 sets all registers to zero on power up.
// Holding reset will set to default values.
reg [7:0] count = 0;
always @ (posedge clk_96mhz)
begin
    if (count < 10) begin
        reset <= 1;
        count <= count + 1;
    end else begin
        reset <= 0;
    end
end

// loopback
reg loop_state;
localparam RECV_CHAR = 0;
localparam SEND_CHAR = 1;
always @ (posedge clk_96mhz)
begin
    if (reset) begin
        uart_rd <= 0;
        uart_wr <= 0;
        tx_data <= 0;
        loop_state <= 0;
        led <= 0;
    end else begin
        case (loop_state)
            RECV_CHAR : begin
                uart_rd <= 0;
                uart_wr <= 0;
                if (rx_valid) begin
                    uart_rd <= 1;
                    tx_data <= rx_data;
                    led <= rx_data;
                    loop_state <= SEND_CHAR;
                end
            end
            SEND_CHAR : begin
                uart_rd <= 0;
                if (~tx_busy) begin
                    uart_wr <= 1;
                    loop_state <= RECV_CHAR;
                end
            end
            default : begin
            end
        endcase
    end
end

endmodule

