// Minimal module
module hello0;
endmodule

