module hello1;
initial $display("Hello World1");
endmodule

