// 0_Input_Output.  Button directly to led.

module top
(
    input wire button0,
    output wire led0
);

assign leds = button0;

endmodule
