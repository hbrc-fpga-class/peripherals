module hello2;
initial 
begin
    $display("Hello World2");
    $display("Goodbye");
end
endmodule

